//Erik Fox
//1/8/2021
//ECE571 - HW1
//Four bit Arbiter (hierarchical/structural)

module Arbiter4(r,g);
input [0:3]r;
output[0:3]g;

endmodule
