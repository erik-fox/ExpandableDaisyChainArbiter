//Erik Fox
//1/8/2021
//ECE571-HW 1
//Four Bit Arbiter, Behavioral model


module Arbiter4(r,g);
input [0:3]r;
input [0:3]g;

endmodule
