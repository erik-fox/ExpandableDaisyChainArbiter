//Erik Fox
//1/8/2021
//ECE571 - HW 1
//Four bit arbiter Testbench

module top;


endmodule
